module CGRA_configurator(
    input      clock,
    input      enable,
    input      sync_reset,

    output reg bitstream,
    output reg done
);

    localparam TOTAL_NUM_BITS = 5821;
	reg [0:TOTAL_NUM_BITS-1] storage = {
		1'bx,1'bx,1'bx, // crossbar::Mux6config
		1'bx,1'bx,1'bx, // crossbar::Mux5config
		1'bx,1'bx,1'bx, // crossbar::Mux4config
		1'bx,1'bx,1'bx, // crossbar::Mux3config
		1'bx,1'bx,1'bx, // crossbar::Mux2config
		1'bx,1'bx,1'bx, // crossbar::Mux1config
		1'bx,1'bx,1'bx, // crossbar::Mux0config
		1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0, // pe_c7_r7::ConstVal
		1'bx, // pe_c7_r7::RegBConfig
		1'bx, // pe_c7_r7::RegAConfig
		1'bx, // pe_c7_r7::Reg4config
		1'bx, // pe_c7_r7::Reg3config
		1'bx, // pe_c7_r7::Reg2config
		1'bx, // pe_c7_r7::Reg1config
		1'bx, // pe_c7_r7::Reg0config
		1'bx, // pe_c7_r7::RESConfig
		1'bx, // pe_c7_r7::Mux4config
		1'bx, // pe_c7_r7::Mux3config
		1'bx, // pe_c7_r7::Mux2config
		1'bx, // pe_c7_r7::Mux1config
		1'bx, // pe_c7_r7::Mux0config
		1'bx,1'bx,1'bx,1'bx, // pe_c7_r7::ALUconfig
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux7config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux6config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux5config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux4config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux3config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux2config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux1config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux0config
		1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0, // pe_c7_r6::ConstVal
		1'bx, // pe_c7_r6::RegBConfig
		1'bx, // pe_c7_r6::RegAConfig
		1'bx, // pe_c7_r6::Reg7config
		1'bx, // pe_c7_r6::Reg4config
		1'bx, // pe_c7_r6::Reg3config
		1'bx, // pe_c7_r6::Reg2config
		1'bx, // pe_c7_r6::Reg1config
		1'bx, // pe_c7_r6::Reg0config
		1'bx, // pe_c7_r6::RESConfig
		1'bx, // pe_c7_r6::Mux7config
		1'bx, // pe_c7_r6::Mux4config
		1'bx, // pe_c7_r6::Mux3config
		1'bx, // pe_c7_r6::Mux2config
		1'bx, // pe_c7_r6::Mux1config
		1'bx, // pe_c7_r6::Mux0config
		1'bx,1'bx,1'bx,1'bx, // pe_c7_r6::ALUconfig
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux7config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux6config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux5config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux4config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux3config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux2config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux1config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux0config
		1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0, // pe_c7_r5::ConstVal
		1'bx, // pe_c7_r5::RegBConfig
		1'bx, // pe_c7_r5::RegAConfig
		1'bx, // pe_c7_r5::Reg7config
		1'bx, // pe_c7_r5::Reg4config
		1'bx, // pe_c7_r5::Reg3config
		1'bx, // pe_c7_r5::Reg2config
		1'bx, // pe_c7_r5::Reg1config
		1'bx, // pe_c7_r5::Reg0config
		1'bx, // pe_c7_r5::RESConfig
		1'bx, // pe_c7_r5::Mux7config
		1'bx, // pe_c7_r5::Mux4config
		1'bx, // pe_c7_r5::Mux3config
		1'bx, // pe_c7_r5::Mux2config
		1'bx, // pe_c7_r5::Mux1config
		1'bx, // pe_c7_r5::Mux0config
		1'bx,1'bx,1'bx,1'bx, // pe_c7_r5::ALUconfig
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux7config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux6config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux5config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux4config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux3config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux2config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux1config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux0config
		1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0, // pe_c7_r4::ConstVal
		1'bx, // pe_c7_r4::RegBConfig
		1'bx, // pe_c7_r4::RegAConfig
		1'bx, // pe_c7_r4::Reg7config
		1'bx, // pe_c7_r4::Reg4config
		1'bx, // pe_c7_r4::Reg3config
		1'bx, // pe_c7_r4::Reg2config
		1'bx, // pe_c7_r4::Reg1config
		1'bx, // pe_c7_r4::Reg0config
		1'bx, // pe_c7_r4::RESConfig
		1'bx, // pe_c7_r4::Mux7config
		1'bx, // pe_c7_r4::Mux4config
		1'bx, // pe_c7_r4::Mux3config
		1'bx, // pe_c7_r4::Mux2config
		1'bx, // pe_c7_r4::Mux1config
		1'bx, // pe_c7_r4::Mux0config
		1'bx,1'bx,1'bx,1'bx, // pe_c7_r4::ALUconfig
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux7config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux6config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux5config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux4config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux3config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux2config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux1config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux0config
		1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0, // pe_c7_r3::ConstVal
		1'bx, // pe_c7_r3::RegBConfig
		1'bx, // pe_c7_r3::RegAConfig
		1'bx, // pe_c7_r3::Reg7config
		1'bx, // pe_c7_r3::Reg4config
		1'bx, // pe_c7_r3::Reg3config
		1'bx, // pe_c7_r3::Reg2config
		1'bx, // pe_c7_r3::Reg1config
		1'bx, // pe_c7_r3::Reg0config
		1'bx, // pe_c7_r3::RESConfig
		1'bx, // pe_c7_r3::Mux7config
		1'bx, // pe_c7_r3::Mux4config
		1'bx, // pe_c7_r3::Mux3config
		1'bx, // pe_c7_r3::Mux2config
		1'bx, // pe_c7_r3::Mux1config
		1'bx, // pe_c7_r3::Mux0config
		1'bx,1'bx,1'bx,1'bx, // pe_c7_r3::ALUconfig
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux7config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux6config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux5config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux4config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux3config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux2config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux1config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux0config
		1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0, // pe_c7_r2::ConstVal
		1'bx, // pe_c7_r2::RegBConfig
		1'bx, // pe_c7_r2::RegAConfig
		1'bx, // pe_c7_r2::Reg7config
		1'bx, // pe_c7_r2::Reg4config
		1'bx, // pe_c7_r2::Reg3config
		1'bx, // pe_c7_r2::Reg2config
		1'bx, // pe_c7_r2::Reg1config
		1'bx, // pe_c7_r2::Reg0config
		1'bx, // pe_c7_r2::RESConfig
		1'bx, // pe_c7_r2::Mux7config
		1'bx, // pe_c7_r2::Mux4config
		1'bx, // pe_c7_r2::Mux3config
		1'bx, // pe_c7_r2::Mux2config
		1'bx, // pe_c7_r2::Mux1config
		1'bx, // pe_c7_r2::Mux0config
		1'bx,1'bx,1'bx,1'bx, // pe_c7_r2::ALUconfig
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux7config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux6config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux5config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux4config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux3config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux2config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux1config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux0config
		1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0, // pe_c7_r1::ConstVal
		1'bx, // pe_c7_r1::RegBConfig
		1'bx, // pe_c7_r1::RegAConfig
		1'bx, // pe_c7_r1::Reg7config
		1'bx, // pe_c7_r1::Reg4config
		1'bx, // pe_c7_r1::Reg3config
		1'bx, // pe_c7_r1::Reg2config
		1'bx, // pe_c7_r1::Reg1config
		1'bx, // pe_c7_r1::Reg0config
		1'bx, // pe_c7_r1::RESConfig
		1'bx, // pe_c7_r1::Mux7config
		1'bx, // pe_c7_r1::Mux4config
		1'bx, // pe_c7_r1::Mux3config
		1'bx, // pe_c7_r1::Mux2config
		1'bx, // pe_c7_r1::Mux1config
		1'bx, // pe_c7_r1::Mux0config
		1'bx,1'bx,1'bx,1'bx, // pe_c7_r1::ALUconfig
		1'bx,1'bx,1'bx, // crossbar::Mux6config
		1'bx,1'bx,1'bx, // crossbar::Mux5config
		1'bx,1'bx,1'bx, // crossbar::Mux4config
		1'b1,1'b1,1'b1, // crossbar::Mux3config
		1'bx,1'bx,1'bx, // crossbar::Mux2config
		1'bx,1'bx,1'bx, // crossbar::Mux1config
		1'bx,1'bx,1'bx, // crossbar::Mux0config
		1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0, // pe_c7_r0::ConstVal
		1'bx, // pe_c7_r0::RegBConfig
		1'bx, // pe_c7_r0::RegAConfig
		1'bx, // pe_c7_r0::Reg7config
		1'bx, // pe_c7_r0::Reg3config
		1'bx, // pe_c7_r0::Reg2config
		1'bx, // pe_c7_r0::Reg1config
		1'bx, // pe_c7_r0::Reg0config
		1'bx, // pe_c7_r0::RESConfig
		1'bx, // pe_c7_r0::Mux7config
		1'bx, // pe_c7_r0::Mux3config
		1'bx, // pe_c7_r0::Mux2config
		1'bx, // pe_c7_r0::Mux1config
		1'bx, // pe_c7_r0::Mux0config
		1'bx,1'bx,1'bx,1'bx, // pe_c7_r0::ALUconfig
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux7config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux6config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux5config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux4config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux3config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux2config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux1config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux0config
		1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0, // pe_c6_r7::ConstVal
		1'bx, // pe_c6_r7::RegBConfig
		1'bx, // pe_c6_r7::RegAConfig
		1'bx, // pe_c6_r7::Reg5config
		1'bx, // pe_c6_r7::Reg4config
		1'bx, // pe_c6_r7::Reg3config
		1'bx, // pe_c6_r7::Reg2config
		1'bx, // pe_c6_r7::Reg1config
		1'bx, // pe_c6_r7::Reg0config
		1'bx, // pe_c6_r7::RESConfig
		1'bx, // pe_c6_r7::Mux5config
		1'bx, // pe_c6_r7::Mux4config
		1'bx, // pe_c6_r7::Mux3config
		1'bx, // pe_c6_r7::Mux2config
		1'bx, // pe_c6_r7::Mux1config
		1'bx, // pe_c6_r7::Mux0config
		1'bx,1'bx,1'bx,1'bx, // pe_c6_r7::ALUconfig
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux9config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux8config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux7config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux6config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux5config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux4config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux3config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux2config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux1config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux0config
		1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0, // pe_c6_r6::ConstVal
		1'bx, // pe_c6_r6::RegBConfig
		1'bx, // pe_c6_r6::RegAConfig
		1'bx, // pe_c6_r6::Reg7config
		1'bx, // pe_c6_r6::Reg6config
		1'bx, // pe_c6_r6::Reg5config
		1'bx, // pe_c6_r6::Reg4config
		1'bx, // pe_c6_r6::Reg3config
		1'bx, // pe_c6_r6::Reg2config
		1'bx, // pe_c6_r6::Reg1config
		1'bx, // pe_c6_r6::Reg0config
		1'bx, // pe_c6_r6::RESConfig
		1'bx, // pe_c6_r6::Mux7config
		1'bx, // pe_c6_r6::Mux6config
		1'bx, // pe_c6_r6::Mux5config
		1'bx, // pe_c6_r6::Mux4config
		1'bx, // pe_c6_r6::Mux3config
		1'bx, // pe_c6_r6::Mux2config
		1'bx, // pe_c6_r6::Mux1config
		1'bx, // pe_c6_r6::Mux0config
		1'bx,1'bx,1'bx,1'bx, // pe_c6_r6::ALUconfig
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux9config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux8config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux7config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux6config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux5config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux4config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux3config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux2config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux1config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux0config
		1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0, // pe_c6_r5::ConstVal
		1'bx, // pe_c6_r5::RegBConfig
		1'bx, // pe_c6_r5::RegAConfig
		1'bx, // pe_c6_r5::Reg7config
		1'bx, // pe_c6_r5::Reg6config
		1'bx, // pe_c6_r5::Reg5config
		1'bx, // pe_c6_r5::Reg4config
		1'bx, // pe_c6_r5::Reg3config
		1'bx, // pe_c6_r5::Reg2config
		1'bx, // pe_c6_r5::Reg1config
		1'bx, // pe_c6_r5::Reg0config
		1'bx, // pe_c6_r5::RESConfig
		1'bx, // pe_c6_r5::Mux7config
		1'bx, // pe_c6_r5::Mux6config
		1'bx, // pe_c6_r5::Mux5config
		1'bx, // pe_c6_r5::Mux4config
		1'bx, // pe_c6_r5::Mux3config
		1'bx, // pe_c6_r5::Mux2config
		1'bx, // pe_c6_r5::Mux1config
		1'bx, // pe_c6_r5::Mux0config
		1'bx,1'bx,1'bx,1'bx, // pe_c6_r5::ALUconfig
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux9config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux8config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux7config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux6config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux5config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux4config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux3config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux2config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux1config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux0config
		1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0, // pe_c6_r4::ConstVal
		1'bx, // pe_c6_r4::RegBConfig
		1'bx, // pe_c6_r4::RegAConfig
		1'bx, // pe_c6_r4::Reg7config
		1'bx, // pe_c6_r4::Reg6config
		1'bx, // pe_c6_r4::Reg5config
		1'bx, // pe_c6_r4::Reg4config
		1'bx, // pe_c6_r4::Reg3config
		1'bx, // pe_c6_r4::Reg2config
		1'bx, // pe_c6_r4::Reg1config
		1'bx, // pe_c6_r4::Reg0config
		1'bx, // pe_c6_r4::RESConfig
		1'bx, // pe_c6_r4::Mux7config
		1'bx, // pe_c6_r4::Mux6config
		1'bx, // pe_c6_r4::Mux5config
		1'bx, // pe_c6_r4::Mux4config
		1'bx, // pe_c6_r4::Mux3config
		1'bx, // pe_c6_r4::Mux2config
		1'bx, // pe_c6_r4::Mux1config
		1'bx, // pe_c6_r4::Mux0config
		1'bx,1'bx,1'bx,1'bx, // pe_c6_r4::ALUconfig
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux9config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux8config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux7config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux6config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux5config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux4config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux3config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux2config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux1config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux0config
		1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0, // pe_c6_r3::ConstVal
		1'bx, // pe_c6_r3::RegBConfig
		1'bx, // pe_c6_r3::RegAConfig
		1'bx, // pe_c6_r3::Reg7config
		1'bx, // pe_c6_r3::Reg6config
		1'bx, // pe_c6_r3::Reg5config
		1'bx, // pe_c6_r3::Reg4config
		1'bx, // pe_c6_r3::Reg3config
		1'bx, // pe_c6_r3::Reg2config
		1'bx, // pe_c6_r3::Reg1config
		1'bx, // pe_c6_r3::Reg0config
		1'bx, // pe_c6_r3::RESConfig
		1'bx, // pe_c6_r3::Mux7config
		1'bx, // pe_c6_r3::Mux6config
		1'bx, // pe_c6_r3::Mux5config
		1'bx, // pe_c6_r3::Mux4config
		1'bx, // pe_c6_r3::Mux3config
		1'bx, // pe_c6_r3::Mux2config
		1'bx, // pe_c6_r3::Mux1config
		1'bx, // pe_c6_r3::Mux0config
		1'bx,1'bx,1'bx,1'bx, // pe_c6_r3::ALUconfig
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux9config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux8config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux7config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux6config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux5config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux4config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux3config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux2config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux1config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux0config
		1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0, // pe_c6_r2::ConstVal
		1'bx, // pe_c6_r2::RegBConfig
		1'bx, // pe_c6_r2::RegAConfig
		1'bx, // pe_c6_r2::Reg7config
		1'bx, // pe_c6_r2::Reg6config
		1'bx, // pe_c6_r2::Reg5config
		1'bx, // pe_c6_r2::Reg4config
		1'bx, // pe_c6_r2::Reg3config
		1'bx, // pe_c6_r2::Reg2config
		1'bx, // pe_c6_r2::Reg1config
		1'bx, // pe_c6_r2::Reg0config
		1'bx, // pe_c6_r2::RESConfig
		1'bx, // pe_c6_r2::Mux7config
		1'bx, // pe_c6_r2::Mux6config
		1'bx, // pe_c6_r2::Mux5config
		1'bx, // pe_c6_r2::Mux4config
		1'bx, // pe_c6_r2::Mux3config
		1'bx, // pe_c6_r2::Mux2config
		1'bx, // pe_c6_r2::Mux1config
		1'bx, // pe_c6_r2::Mux0config
		1'bx,1'bx,1'bx,1'bx, // pe_c6_r2::ALUconfig
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux9config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux8config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux7config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux6config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux5config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux4config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux3config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux2config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux1config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux0config
		1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0, // pe_c6_r1::ConstVal
		1'bx, // pe_c6_r1::RegBConfig
		1'bx, // pe_c6_r1::RegAConfig
		1'bx, // pe_c6_r1::Reg7config
		1'bx, // pe_c6_r1::Reg6config
		1'bx, // pe_c6_r1::Reg5config
		1'bx, // pe_c6_r1::Reg4config
		1'bx, // pe_c6_r1::Reg3config
		1'bx, // pe_c6_r1::Reg2config
		1'bx, // pe_c6_r1::Reg1config
		1'bx, // pe_c6_r1::Reg0config
		1'bx, // pe_c6_r1::RESConfig
		1'bx, // pe_c6_r1::Mux7config
		1'bx, // pe_c6_r1::Mux6config
		1'bx, // pe_c6_r1::Mux5config
		1'bx, // pe_c6_r1::Mux4config
		1'bx, // pe_c6_r1::Mux3config
		1'bx, // pe_c6_r1::Mux2config
		1'bx, // pe_c6_r1::Mux1config
		1'bx, // pe_c6_r1::Mux0config
		1'bx,1'bx,1'bx,1'bx, // pe_c6_r1::ALUconfig
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux7config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux6config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux5config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux4config
		1'b1,1'b0,1'b0,1'b0, // crossbar::Mux3config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux2config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux1config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux0config
		1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0, // pe_c6_r0::ConstVal
		1'bx, // pe_c6_r0::RegBConfig
		1'bx, // pe_c6_r0::RegAConfig
		1'bx, // pe_c6_r0::Reg7config
		1'bx, // pe_c6_r0::Reg6config
		1'bx, // pe_c6_r0::Reg3config
		1'bx, // pe_c6_r0::Reg2config
		1'bx, // pe_c6_r0::Reg1config
		1'bx, // pe_c6_r0::Reg0config
		1'bx, // pe_c6_r0::RESConfig
		1'bx, // pe_c6_r0::Mux7config
		1'bx, // pe_c6_r0::Mux6config
		1'bx, // pe_c6_r0::Mux3config
		1'bx, // pe_c6_r0::Mux2config
		1'b0, // pe_c6_r0::Mux1config
		1'bx, // pe_c6_r0::Mux0config
		1'bx,1'bx,1'bx,1'bx, // pe_c6_r0::ALUconfig
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux7config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux6config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux5config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux4config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux3config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux2config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux1config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux0config
		1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0, // pe_c5_r7::ConstVal
		1'bx, // pe_c5_r7::RegBConfig
		1'bx, // pe_c5_r7::RegAConfig
		1'bx, // pe_c5_r7::Reg5config
		1'bx, // pe_c5_r7::Reg4config
		1'bx, // pe_c5_r7::Reg3config
		1'bx, // pe_c5_r7::Reg2config
		1'bx, // pe_c5_r7::Reg1config
		1'bx, // pe_c5_r7::Reg0config
		1'bx, // pe_c5_r7::RESConfig
		1'bx, // pe_c5_r7::Mux5config
		1'bx, // pe_c5_r7::Mux4config
		1'bx, // pe_c5_r7::Mux3config
		1'bx, // pe_c5_r7::Mux2config
		1'bx, // pe_c5_r7::Mux1config
		1'bx, // pe_c5_r7::Mux0config
		1'bx,1'bx,1'bx,1'bx, // pe_c5_r7::ALUconfig
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux9config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux8config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux7config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux6config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux5config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux4config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux3config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux2config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux1config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux0config
		1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0, // pe_c5_r6::ConstVal
		1'bx, // pe_c5_r6::RegBConfig
		1'bx, // pe_c5_r6::RegAConfig
		1'bx, // pe_c5_r6::Reg7config
		1'bx, // pe_c5_r6::Reg6config
		1'bx, // pe_c5_r6::Reg5config
		1'bx, // pe_c5_r6::Reg4config
		1'bx, // pe_c5_r6::Reg3config
		1'bx, // pe_c5_r6::Reg2config
		1'bx, // pe_c5_r6::Reg1config
		1'bx, // pe_c5_r6::Reg0config
		1'bx, // pe_c5_r6::RESConfig
		1'bx, // pe_c5_r6::Mux7config
		1'bx, // pe_c5_r6::Mux6config
		1'bx, // pe_c5_r6::Mux5config
		1'bx, // pe_c5_r6::Mux4config
		1'bx, // pe_c5_r6::Mux3config
		1'bx, // pe_c5_r6::Mux2config
		1'bx, // pe_c5_r6::Mux1config
		1'bx, // pe_c5_r6::Mux0config
		1'bx,1'bx,1'bx,1'bx, // pe_c5_r6::ALUconfig
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux9config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux8config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux7config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux6config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux5config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux4config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux3config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux2config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux1config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux0config
		1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0, // pe_c5_r5::ConstVal
		1'bx, // pe_c5_r5::RegBConfig
		1'bx, // pe_c5_r5::RegAConfig
		1'bx, // pe_c5_r5::Reg7config
		1'bx, // pe_c5_r5::Reg6config
		1'bx, // pe_c5_r5::Reg5config
		1'bx, // pe_c5_r5::Reg4config
		1'bx, // pe_c5_r5::Reg3config
		1'bx, // pe_c5_r5::Reg2config
		1'bx, // pe_c5_r5::Reg1config
		1'bx, // pe_c5_r5::Reg0config
		1'bx, // pe_c5_r5::RESConfig
		1'bx, // pe_c5_r5::Mux7config
		1'bx, // pe_c5_r5::Mux6config
		1'bx, // pe_c5_r5::Mux5config
		1'bx, // pe_c5_r5::Mux4config
		1'bx, // pe_c5_r5::Mux3config
		1'bx, // pe_c5_r5::Mux2config
		1'bx, // pe_c5_r5::Mux1config
		1'bx, // pe_c5_r5::Mux0config
		1'bx,1'bx,1'bx,1'bx, // pe_c5_r5::ALUconfig
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux9config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux8config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux7config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux6config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux5config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux4config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux3config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux2config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux1config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux0config
		1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0, // pe_c5_r4::ConstVal
		1'bx, // pe_c5_r4::RegBConfig
		1'bx, // pe_c5_r4::RegAConfig
		1'bx, // pe_c5_r4::Reg7config
		1'bx, // pe_c5_r4::Reg6config
		1'bx, // pe_c5_r4::Reg5config
		1'bx, // pe_c5_r4::Reg4config
		1'bx, // pe_c5_r4::Reg3config
		1'bx, // pe_c5_r4::Reg2config
		1'bx, // pe_c5_r4::Reg1config
		1'bx, // pe_c5_r4::Reg0config
		1'bx, // pe_c5_r4::RESConfig
		1'bx, // pe_c5_r4::Mux7config
		1'bx, // pe_c5_r4::Mux6config
		1'bx, // pe_c5_r4::Mux5config
		1'bx, // pe_c5_r4::Mux4config
		1'bx, // pe_c5_r4::Mux3config
		1'bx, // pe_c5_r4::Mux2config
		1'bx, // pe_c5_r4::Mux1config
		1'bx, // pe_c5_r4::Mux0config
		1'bx,1'bx,1'bx,1'bx, // pe_c5_r4::ALUconfig
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux9config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux8config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux7config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux6config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux5config
		1'b0,1'b1,1'b0,1'b1, // crossbar::Mux4config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux3config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux2config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux1config
		1'b1,1'b1,1'b0,1'b0, // crossbar::Mux0config
		1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0, // pe_c5_r3::ConstVal
		1'bx, // pe_c5_r3::RegBConfig
		1'bx, // pe_c5_r3::RegAConfig
		1'bx, // pe_c5_r3::Reg7config
		1'bx, // pe_c5_r3::Reg6config
		1'bx, // pe_c5_r3::Reg5config
		1'bx, // pe_c5_r3::Reg4config
		1'bx, // pe_c5_r3::Reg3config
		1'bx, // pe_c5_r3::Reg2config
		1'bx, // pe_c5_r3::Reg1config
		1'bx, // pe_c5_r3::Reg0config
		1'bx, // pe_c5_r3::RESConfig
		1'bx, // pe_c5_r3::Mux7config
		1'bx, // pe_c5_r3::Mux6config
		1'bx, // pe_c5_r3::Mux5config
		1'bx, // pe_c5_r3::Mux4config
		1'b0, // pe_c5_r3::Mux3config
		1'bx, // pe_c5_r3::Mux2config
		1'bx, // pe_c5_r3::Mux1config
		1'bx, // pe_c5_r3::Mux0config
		1'bx,1'bx,1'bx,1'bx, // pe_c5_r3::ALUconfig
		1'b0,1'b1,1'b0,1'b0, // crossbar::Mux9config
		1'b1,1'b1,1'b1,1'b0, // crossbar::Mux8config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux7config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux6config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux5config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux4config
		1'b0,1'b0,1'b0,1'b1, // crossbar::Mux3config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux2config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux1config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux0config
		1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0, // pe_c5_r2::ConstVal
		1'b1, // pe_c5_r2::RegBConfig
		1'b1, // pe_c5_r2::RegAConfig
		1'bx, // pe_c5_r2::Reg7config
		1'bx, // pe_c5_r2::Reg6config
		1'bx, // pe_c5_r2::Reg5config
		1'bx, // pe_c5_r2::Reg4config
		1'bx, // pe_c5_r2::Reg3config
		1'bx, // pe_c5_r2::Reg2config
		1'bx, // pe_c5_r2::Reg1config
		1'bx, // pe_c5_r2::Reg0config
		1'bx, // pe_c5_r2::RESConfig
		1'b0, // pe_c5_r2::Mux7config
		1'bx, // pe_c5_r2::Mux6config
		1'bx, // pe_c5_r2::Mux5config
		1'bx, // pe_c5_r2::Mux4config
		1'bx, // pe_c5_r2::Mux3config
		1'b0, // pe_c5_r2::Mux2config
		1'bx, // pe_c5_r2::Mux1config
		1'bx, // pe_c5_r2::Mux0config
		1'b0,1'b0,1'b0,1'b0, // pe_c5_r2::ALUconfig
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux9config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux8config
		1'b0,1'b0,1'b0,1'b0, // crossbar::Mux7config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux6config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux5config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux4config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux3config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux2config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux1config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux0config
		1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0, // pe_c5_r1::ConstVal
		1'bx, // pe_c5_r1::RegBConfig
		1'bx, // pe_c5_r1::RegAConfig
		1'bx, // pe_c5_r1::Reg7config
		1'bx, // pe_c5_r1::Reg6config
		1'bx, // pe_c5_r1::Reg5config
		1'bx, // pe_c5_r1::Reg4config
		1'bx, // pe_c5_r1::Reg3config
		1'bx, // pe_c5_r1::Reg2config
		1'bx, // pe_c5_r1::Reg1config
		1'bx, // pe_c5_r1::Reg0config
		1'bx, // pe_c5_r1::RESConfig
		1'bx, // pe_c5_r1::Mux7config
		1'bx, // pe_c5_r1::Mux6config
		1'bx, // pe_c5_r1::Mux5config
		1'bx, // pe_c5_r1::Mux4config
		1'bx, // pe_c5_r1::Mux3config
		1'bx, // pe_c5_r1::Mux2config
		1'bx, // pe_c5_r1::Mux1config
		1'b0, // pe_c5_r1::Mux0config
		1'bx,1'bx,1'bx,1'bx, // pe_c5_r1::ALUconfig
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux7config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux6config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux5config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux4config
		1'b1,1'b0,1'b0,1'b0, // crossbar::Mux3config
		1'b0,1'b0,1'b0,1'b1, // crossbar::Mux2config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux1config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux0config
		1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0, // pe_c5_r0::ConstVal
		1'bx, // pe_c5_r0::RegBConfig
		1'bx, // pe_c5_r0::RegAConfig
		1'bx, // pe_c5_r0::Reg7config
		1'bx, // pe_c5_r0::Reg6config
		1'bx, // pe_c5_r0::Reg3config
		1'bx, // pe_c5_r0::Reg2config
		1'bx, // pe_c5_r0::Reg1config
		1'bx, // pe_c5_r0::Reg0config
		1'bx, // pe_c5_r0::RESConfig
		1'bx, // pe_c5_r0::Mux7config
		1'bx, // pe_c5_r0::Mux6config
		1'bx, // pe_c5_r0::Mux3config
		1'bx, // pe_c5_r0::Mux2config
		1'b0, // pe_c5_r0::Mux1config
		1'bx, // pe_c5_r0::Mux0config
		1'bx,1'bx,1'bx,1'bx, // pe_c5_r0::ALUconfig
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux7config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux6config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux5config
		1'b0,1'b0,1'b0,1'b0, // crossbar::Mux4config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux3config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux2config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux1config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux0config
		1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0, // pe_c4_r7::ConstVal
		1'bx, // pe_c4_r7::RegBConfig
		1'bx, // pe_c4_r7::RegAConfig
		1'bx, // pe_c4_r7::Reg5config
		1'bx, // pe_c4_r7::Reg4config
		1'bx, // pe_c4_r7::Reg3config
		1'bx, // pe_c4_r7::Reg2config
		1'bx, // pe_c4_r7::Reg1config
		1'bx, // pe_c4_r7::Reg0config
		1'bx, // pe_c4_r7::RESConfig
		1'bx, // pe_c4_r7::Mux5config
		1'bx, // pe_c4_r7::Mux4config
		1'bx, // pe_c4_r7::Mux3config
		1'bx, // pe_c4_r7::Mux2config
		1'bx, // pe_c4_r7::Mux1config
		1'b0, // pe_c4_r7::Mux0config
		1'bx,1'bx,1'bx,1'bx, // pe_c4_r7::ALUconfig
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux9config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux8config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux7config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux6config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux5config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux4config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux3config
		1'b0,1'b1,1'b0,1'b1, // crossbar::Mux2config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux1config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux0config
		1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0, // pe_c4_r6::ConstVal
		1'bx, // pe_c4_r6::RegBConfig
		1'bx, // pe_c4_r6::RegAConfig
		1'bx, // pe_c4_r6::Reg7config
		1'bx, // pe_c4_r6::Reg6config
		1'bx, // pe_c4_r6::Reg5config
		1'bx, // pe_c4_r6::Reg4config
		1'bx, // pe_c4_r6::Reg3config
		1'bx, // pe_c4_r6::Reg2config
		1'bx, // pe_c4_r6::Reg1config
		1'bx, // pe_c4_r6::Reg0config
		1'bx, // pe_c4_r6::RESConfig
		1'bx, // pe_c4_r6::Mux7config
		1'bx, // pe_c4_r6::Mux6config
		1'bx, // pe_c4_r6::Mux5config
		1'bx, // pe_c4_r6::Mux4config
		1'bx, // pe_c4_r6::Mux3config
		1'bx, // pe_c4_r6::Mux2config
		1'bx, // pe_c4_r6::Mux1config
		1'bx, // pe_c4_r6::Mux0config
		1'bx,1'bx,1'bx,1'bx, // pe_c4_r6::ALUconfig
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux9config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux8config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux7config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux6config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux5config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux4config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux3config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux2config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux1config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux0config
		1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0, // pe_c4_r5::ConstVal
		1'bx, // pe_c4_r5::RegBConfig
		1'bx, // pe_c4_r5::RegAConfig
		1'bx, // pe_c4_r5::Reg7config
		1'bx, // pe_c4_r5::Reg6config
		1'bx, // pe_c4_r5::Reg5config
		1'bx, // pe_c4_r5::Reg4config
		1'bx, // pe_c4_r5::Reg3config
		1'bx, // pe_c4_r5::Reg2config
		1'bx, // pe_c4_r5::Reg1config
		1'bx, // pe_c4_r5::Reg0config
		1'bx, // pe_c4_r5::RESConfig
		1'bx, // pe_c4_r5::Mux7config
		1'bx, // pe_c4_r5::Mux6config
		1'bx, // pe_c4_r5::Mux5config
		1'bx, // pe_c4_r5::Mux4config
		1'bx, // pe_c4_r5::Mux3config
		1'bx, // pe_c4_r5::Mux2config
		1'bx, // pe_c4_r5::Mux1config
		1'bx, // pe_c4_r5::Mux0config
		1'bx,1'bx,1'bx,1'bx, // pe_c4_r5::ALUconfig
		1'b0,1'b0,1'b1,1'b0, // crossbar::Mux9config
		1'b1,1'b1,1'b0,1'b0, // crossbar::Mux8config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux7config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux6config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux5config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux4config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux3config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux2config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux1config
		1'b0,1'b0,1'b0,1'b1, // crossbar::Mux0config
		1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0, // pe_c4_r4::ConstVal
		1'b1, // pe_c4_r4::RegBConfig
		1'b1, // pe_c4_r4::RegAConfig
		1'bx, // pe_c4_r4::Reg7config
		1'bx, // pe_c4_r4::Reg6config
		1'bx, // pe_c4_r4::Reg5config
		1'bx, // pe_c4_r4::Reg4config
		1'bx, // pe_c4_r4::Reg3config
		1'bx, // pe_c4_r4::Reg2config
		1'bx, // pe_c4_r4::Reg1config
		1'bx, // pe_c4_r4::Reg0config
		1'bx, // pe_c4_r4::RESConfig
		1'bx, // pe_c4_r4::Mux7config
		1'bx, // pe_c4_r4::Mux6config
		1'bx, // pe_c4_r4::Mux5config
		1'b0, // pe_c4_r4::Mux4config
		1'b0, // pe_c4_r4::Mux3config
		1'bx, // pe_c4_r4::Mux2config
		1'bx, // pe_c4_r4::Mux1config
		1'bx, // pe_c4_r4::Mux0config
		1'b0,1'b1,1'b0,1'b0, // pe_c4_r4::ALUconfig
		1'b1,1'b1,1'b1,1'b0, // crossbar::Mux9config
		1'b0,1'b0,1'b1,1'b0, // crossbar::Mux8config
		1'b1,1'b1,1'b0,1'b0, // crossbar::Mux7config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux6config
		1'b0,1'b1,1'b0,1'b0, // crossbar::Mux5config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux4config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux3config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux2config
		1'b0,1'b0,1'b0,1'b1, // crossbar::Mux1config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux0config
		1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0, // pe_c4_r3::ConstVal
		1'b1, // pe_c4_r3::RegBConfig
		1'b1, // pe_c4_r3::RegAConfig
		1'bx, // pe_c4_r3::Reg7config
		1'bx, // pe_c4_r3::Reg6config
		1'bx, // pe_c4_r3::Reg5config
		1'b1, // pe_c4_r3::Reg4config
		1'bx, // pe_c4_r3::Reg3config
		1'b1, // pe_c4_r3::Reg2config
		1'bx, // pe_c4_r3::Reg1config
		1'bx, // pe_c4_r3::Reg0config
		1'bx, // pe_c4_r3::RESConfig
		1'b0, // pe_c4_r3::Mux7config
		1'bx, // pe_c4_r3::Mux6config
		1'bx, // pe_c4_r3::Mux5config
		1'b1, // pe_c4_r3::Mux4config
		1'b0, // pe_c4_r3::Mux3config
		1'b1, // pe_c4_r3::Mux2config
		1'bx, // pe_c4_r3::Mux1config
		1'bx, // pe_c4_r3::Mux0config
		1'b0,1'b1,1'b0,1'b0, // pe_c4_r3::ALUconfig
		1'b0,1'b1,1'b1,1'b0, // crossbar::Mux9config
		1'b1,1'b0,1'b0,1'b0, // crossbar::Mux8config
		1'b1,1'b0,1'b1,1'b0, // crossbar::Mux7config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux6config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux5config
		1'b1,1'b0,1'b0,1'b1, // crossbar::Mux4config
		1'b0,1'b0,1'b0,1'b1, // crossbar::Mux3config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux2config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux1config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux0config
		1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0, // pe_c4_r2::ConstVal
		1'b1, // pe_c4_r2::RegBConfig
		1'b1, // pe_c4_r2::RegAConfig
		1'bx, // pe_c4_r2::Reg7config
		1'b1, // pe_c4_r2::Reg6config
		1'bx, // pe_c4_r2::Reg5config
		1'bx, // pe_c4_r2::Reg4config
		1'bx, // pe_c4_r2::Reg3config
		1'bx, // pe_c4_r2::Reg2config
		1'b1, // pe_c4_r2::Reg1config
		1'bx, // pe_c4_r2::Reg0config
		1'b1, // pe_c4_r2::RESConfig
		1'bx, // pe_c4_r2::Mux7config
		1'b1, // pe_c4_r2::Mux6config
		1'b0, // pe_c4_r2::Mux5config
		1'bx, // pe_c4_r2::Mux4config
		1'bx, // pe_c4_r2::Mux3config
		1'bx, // pe_c4_r2::Mux2config
		1'b1, // pe_c4_r2::Mux1config
		1'bx, // pe_c4_r2::Mux0config
		1'b1,1'b1,1'b1,1'b0, // pe_c4_r2::ALUconfig
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux9config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux8config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux7config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux6config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux5config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux4config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux3config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux2config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux1config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux0config
		1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0, // pe_c4_r1::ConstVal
		1'bx, // pe_c4_r1::RegBConfig
		1'bx, // pe_c4_r1::RegAConfig
		1'bx, // pe_c4_r1::Reg7config
		1'bx, // pe_c4_r1::Reg6config
		1'bx, // pe_c4_r1::Reg5config
		1'bx, // pe_c4_r1::Reg4config
		1'bx, // pe_c4_r1::Reg3config
		1'bx, // pe_c4_r1::Reg2config
		1'bx, // pe_c4_r1::Reg1config
		1'bx, // pe_c4_r1::Reg0config
		1'bx, // pe_c4_r1::RESConfig
		1'bx, // pe_c4_r1::Mux7config
		1'bx, // pe_c4_r1::Mux6config
		1'bx, // pe_c4_r1::Mux5config
		1'bx, // pe_c4_r1::Mux4config
		1'bx, // pe_c4_r1::Mux3config
		1'bx, // pe_c4_r1::Mux2config
		1'bx, // pe_c4_r1::Mux1config
		1'bx, // pe_c4_r1::Mux0config
		1'bx,1'bx,1'bx,1'bx, // pe_c4_r1::ALUconfig
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux7config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux6config
		1'b1,1'b0,1'b0,1'b0, // crossbar::Mux5config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux4config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux3config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux2config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux1config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux0config
		1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0, // pe_c4_r0::ConstVal
		1'bx, // pe_c4_r0::RegBConfig
		1'bx, // pe_c4_r0::RegAConfig
		1'bx, // pe_c4_r0::Reg7config
		1'bx, // pe_c4_r0::Reg6config
		1'bx, // pe_c4_r0::Reg3config
		1'bx, // pe_c4_r0::Reg2config
		1'bx, // pe_c4_r0::Reg1config
		1'bx, // pe_c4_r0::Reg0config
		1'bx, // pe_c4_r0::RESConfig
		1'bx, // pe_c4_r0::Mux7config
		1'bx, // pe_c4_r0::Mux6config
		1'bx, // pe_c4_r0::Mux3config
		1'bx, // pe_c4_r0::Mux2config
		1'b0, // pe_c4_r0::Mux1config
		1'bx, // pe_c4_r0::Mux0config
		1'bx,1'bx,1'bx,1'bx, // pe_c4_r0::ALUconfig
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux7config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux6config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux5config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux4config
		1'b0,1'b1,1'b0,1'b0, // crossbar::Mux3config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux2config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux1config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux0config
		1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0, // pe_c3_r7::ConstVal
		1'bx, // pe_c3_r7::RegBConfig
		1'bx, // pe_c3_r7::RegAConfig
		1'bx, // pe_c3_r7::Reg5config
		1'bx, // pe_c3_r7::Reg4config
		1'bx, // pe_c3_r7::Reg3config
		1'bx, // pe_c3_r7::Reg2config
		1'bx, // pe_c3_r7::Reg1config
		1'bx, // pe_c3_r7::Reg0config
		1'bx, // pe_c3_r7::RESConfig
		1'bx, // pe_c3_r7::Mux5config
		1'bx, // pe_c3_r7::Mux4config
		1'bx, // pe_c3_r7::Mux3config
		1'b0, // pe_c3_r7::Mux2config
		1'bx, // pe_c3_r7::Mux1config
		1'bx, // pe_c3_r7::Mux0config
		1'bx,1'bx,1'bx,1'bx, // pe_c3_r7::ALUconfig
		1'b0,1'b1,1'b1,1'b0, // crossbar::Mux9config
		1'b0,1'b0,1'b1,1'b0, // crossbar::Mux8config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux7config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux6config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux5config
		1'b1,1'b0,1'b0,1'b1, // crossbar::Mux4config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux3config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux2config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux1config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux0config
		1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0, // pe_c3_r6::ConstVal
		1'b1, // pe_c3_r6::RegBConfig
		1'b1, // pe_c3_r6::RegAConfig
		1'bx, // pe_c3_r6::Reg7config
		1'bx, // pe_c3_r6::Reg6config
		1'bx, // pe_c3_r6::Reg5config
		1'bx, // pe_c3_r6::Reg4config
		1'bx, // pe_c3_r6::Reg3config
		1'bx, // pe_c3_r6::Reg2config
		1'bx, // pe_c3_r6::Reg1config
		1'bx, // pe_c3_r6::Reg0config
		1'b1, // pe_c3_r6::RESConfig
		1'bx, // pe_c3_r6::Mux7config
		1'b0, // pe_c3_r6::Mux6config
		1'bx, // pe_c3_r6::Mux5config
		1'b0, // pe_c3_r6::Mux4config
		1'bx, // pe_c3_r6::Mux3config
		1'bx, // pe_c3_r6::Mux2config
		1'bx, // pe_c3_r6::Mux1config
		1'bx, // pe_c3_r6::Mux0config
		1'b1,1'b1,1'b1,1'b0, // pe_c3_r6::ALUconfig
		1'b1,1'b1,1'b1,1'b0, // crossbar::Mux9config
		1'b0,1'b0,1'b1,1'b0, // crossbar::Mux8config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux7config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux6config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux5config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux4config
		1'b1,1'b0,1'b0,1'b1, // crossbar::Mux3config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux2config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux1config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux0config
		1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0, // pe_c3_r5::ConstVal
		1'b1, // pe_c3_r5::RegBConfig
		1'b1, // pe_c3_r5::RegAConfig
		1'b1, // pe_c3_r5::Reg7config
		1'bx, // pe_c3_r5::Reg6config
		1'bx, // pe_c3_r5::Reg5config
		1'bx, // pe_c3_r5::Reg4config
		1'bx, // pe_c3_r5::Reg3config
		1'bx, // pe_c3_r5::Reg2config
		1'bx, // pe_c3_r5::Reg1config
		1'bx, // pe_c3_r5::Reg0config
		1'b1, // pe_c3_r5::RESConfig
		1'b1, // pe_c3_r5::Mux7config
		1'bx, // pe_c3_r5::Mux6config
		1'bx, // pe_c3_r5::Mux5config
		1'b0, // pe_c3_r5::Mux4config
		1'bx, // pe_c3_r5::Mux3config
		1'bx, // pe_c3_r5::Mux2config
		1'bx, // pe_c3_r5::Mux1config
		1'bx, // pe_c3_r5::Mux0config
		1'b0,1'b0,1'b0,1'b1, // pe_c3_r5::ALUconfig
		1'b1,1'b0,1'b1,1'b0, // crossbar::Mux9config
		1'b0,1'b0,1'b0,1'b0, // crossbar::Mux8config
		1'b1,1'b0,1'b0,1'b1, // crossbar::Mux7config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux6config
		1'b1,1'b1,1'b0,1'b0, // crossbar::Mux5config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux4config
		1'b0,1'b1,1'b0,1'b1, // crossbar::Mux3config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux2config
		1'b1,1'b1,1'b1,1'b0, // crossbar::Mux1config
		1'b1,1'b1,1'b1,1'b0, // crossbar::Mux0config
		1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0, // pe_c3_r4::ConstVal
		1'b1, // pe_c3_r4::RegBConfig
		1'b1, // pe_c3_r4::RegAConfig
		1'bx, // pe_c3_r4::Reg7config
		1'bx, // pe_c3_r4::Reg6config
		1'bx, // pe_c3_r4::Reg5config
		1'bx, // pe_c3_r4::Reg4config
		1'b1, // pe_c3_r4::Reg3config
		1'bx, // pe_c3_r4::Reg2config
		1'bx, // pe_c3_r4::Reg1config
		1'bx, // pe_c3_r4::Reg0config
		1'b1, // pe_c3_r4::RESConfig
		1'b0, // pe_c3_r4::Mux7config
		1'bx, // pe_c3_r4::Mux6config
		1'b0, // pe_c3_r4::Mux5config
		1'bx, // pe_c3_r4::Mux4config
		1'b1, // pe_c3_r4::Mux3config
		1'bx, // pe_c3_r4::Mux2config
		1'bx, // pe_c3_r4::Mux1config
		1'b0, // pe_c3_r4::Mux0config
		1'b1,1'b0,1'b0,1'b0, // pe_c3_r4::ALUconfig
		1'b0,1'b1,1'b0,1'b0, // crossbar::Mux9config
		1'b1,1'b1,1'b1,1'b0, // crossbar::Mux8config
		1'b1,1'b0,1'b1,1'b0, // crossbar::Mux7config
		1'b0,1'b0,1'b1,1'b0, // crossbar::Mux6config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux5config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux4config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux3config
		1'b0,1'b0,1'b0,1'b0, // crossbar::Mux2config
		1'b0,1'b0,1'b0,1'b1, // crossbar::Mux1config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux0config
		1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0, // pe_c3_r3::ConstVal
		1'b1, // pe_c3_r3::RegBConfig
		1'b1, // pe_c3_r3::RegAConfig
		1'bx, // pe_c3_r3::Reg7config
		1'bx, // pe_c3_r3::Reg6config
		1'bx, // pe_c3_r3::Reg5config
		1'bx, // pe_c3_r3::Reg4config
		1'bx, // pe_c3_r3::Reg3config
		1'bx, // pe_c3_r3::Reg2config
		1'bx, // pe_c3_r3::Reg1config
		1'bx, // pe_c3_r3::Reg0config
		1'bx, // pe_c3_r3::RESConfig
		1'b0, // pe_c3_r3::Mux7config
		1'bx, // pe_c3_r3::Mux6config
		1'b0, // pe_c3_r3::Mux5config
		1'b0, // pe_c3_r3::Mux4config
		1'bx, // pe_c3_r3::Mux3config
		1'b0, // pe_c3_r3::Mux2config
		1'bx, // pe_c3_r3::Mux1config
		1'b0, // pe_c3_r3::Mux0config
		1'b0,1'b1,1'b0,1'b0, // pe_c3_r3::ALUconfig
		1'b0,1'b0,1'b1,1'b0, // crossbar::Mux9config
		1'b0,1'b0,1'b0,1'b0, // crossbar::Mux8config
		1'b1,1'b0,1'b0,1'b0, // crossbar::Mux7config
		1'b0,1'b0,1'b1,1'b0, // crossbar::Mux6config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux5config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux4config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux3config
		1'b0,1'b0,1'b0,1'b1, // crossbar::Mux2config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux1config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux0config
		1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0, // pe_c3_r2::ConstVal
		1'b1, // pe_c3_r2::RegBConfig
		1'b1, // pe_c3_r2::RegAConfig
		1'bx, // pe_c3_r2::Reg7config
		1'bx, // pe_c3_r2::Reg6config
		1'bx, // pe_c3_r2::Reg5config
		1'bx, // pe_c3_r2::Reg4config
		1'bx, // pe_c3_r2::Reg3config
		1'bx, // pe_c3_r2::Reg2config
		1'bx, // pe_c3_r2::Reg1config
		1'bx, // pe_c3_r2::Reg0config
		1'bx, // pe_c3_r2::RESConfig
		1'bx, // pe_c3_r2::Mux7config
		1'bx, // pe_c3_r2::Mux6config
		1'bx, // pe_c3_r2::Mux5config
		1'b0, // pe_c3_r2::Mux4config
		1'bx, // pe_c3_r2::Mux3config
		1'bx, // pe_c3_r2::Mux2config
		1'b0, // pe_c3_r2::Mux1config
		1'b0, // pe_c3_r2::Mux0config
		1'b0,1'b1,1'b0,1'b0, // pe_c3_r2::ALUconfig
		1'b0,1'b0,1'b1,1'b0, // crossbar::Mux9config
		1'b0,1'b0,1'b0,1'b0, // crossbar::Mux8config
		1'b1,1'b0,1'b1,1'b0, // crossbar::Mux7config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux6config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux5config
		1'b0,1'b1,1'b1,1'b0, // crossbar::Mux4config
		1'b0,1'b0,1'b0,1'b1, // crossbar::Mux3config
		1'b1,1'b1,1'b1,1'b0, // crossbar::Mux2config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux1config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux0config
		1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0, // pe_c3_r1::ConstVal
		1'b1, // pe_c3_r1::RegBConfig
		1'b1, // pe_c3_r1::RegAConfig
		1'bx, // pe_c3_r1::Reg7config
		1'bx, // pe_c3_r1::Reg6config
		1'bx, // pe_c3_r1::Reg5config
		1'b1, // pe_c3_r1::Reg4config
		1'bx, // pe_c3_r1::Reg3config
		1'bx, // pe_c3_r1::Reg2config
		1'bx, // pe_c3_r1::Reg1config
		1'bx, // pe_c3_r1::Reg0config
		1'bx, // pe_c3_r1::RESConfig
		1'b0, // pe_c3_r1::Mux7config
		1'b0, // pe_c3_r1::Mux6config
		1'b0, // pe_c3_r1::Mux5config
		1'b1, // pe_c3_r1::Mux4config
		1'bx, // pe_c3_r1::Mux3config
		1'bx, // pe_c3_r1::Mux2config
		1'bx, // pe_c3_r1::Mux1config
		1'b0, // pe_c3_r1::Mux0config
		1'b0,1'b0,1'b0,1'b1, // pe_c3_r1::ALUconfig
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux7config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux6config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux5config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux4config
		1'b0,1'b0,1'b0,1'b0, // crossbar::Mux3config
		1'b1,1'b1,1'b0,1'b0, // crossbar::Mux2config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux1config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux0config
		1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0, // pe_c3_r0::ConstVal
		1'bx, // pe_c3_r0::RegBConfig
		1'bx, // pe_c3_r0::RegAConfig
		1'bx, // pe_c3_r0::Reg7config
		1'bx, // pe_c3_r0::Reg6config
		1'b1, // pe_c3_r0::Reg3config
		1'bx, // pe_c3_r0::Reg2config
		1'bx, // pe_c3_r0::Reg1config
		1'bx, // pe_c3_r0::Reg0config
		1'bx, // pe_c3_r0::RESConfig
		1'bx, // pe_c3_r0::Mux7config
		1'bx, // pe_c3_r0::Mux6config
		1'b1, // pe_c3_r0::Mux3config
		1'bx, // pe_c3_r0::Mux2config
		1'bx, // pe_c3_r0::Mux1config
		1'b0, // pe_c3_r0::Mux0config
		1'bx,1'bx,1'bx,1'bx, // pe_c3_r0::ALUconfig
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux7config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux6config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux5config
		1'b0,1'b0,1'b0,1'b1, // crossbar::Mux4config
		1'b1,1'b0,1'b0,1'b0, // crossbar::Mux3config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux2config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux1config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux0config
		1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0, // pe_c2_r7::ConstVal
		1'bx, // pe_c2_r7::RegBConfig
		1'bx, // pe_c2_r7::RegAConfig
		1'bx, // pe_c2_r7::Reg5config
		1'bx, // pe_c2_r7::Reg4config
		1'bx, // pe_c2_r7::Reg3config
		1'bx, // pe_c2_r7::Reg2config
		1'bx, // pe_c2_r7::Reg1config
		1'bx, // pe_c2_r7::Reg0config
		1'bx, // pe_c2_r7::RESConfig
		1'bx, // pe_c2_r7::Mux5config
		1'bx, // pe_c2_r7::Mux4config
		1'bx, // pe_c2_r7::Mux3config
		1'bx, // pe_c2_r7::Mux2config
		1'b0, // pe_c2_r7::Mux1config
		1'bx, // pe_c2_r7::Mux0config
		1'bx,1'bx,1'bx,1'bx, // pe_c2_r7::ALUconfig
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux9config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux8config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux7config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux6config
		1'b1,1'b1,1'b1,1'b0, // crossbar::Mux5config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux4config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux3config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux2config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux1config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux0config
		1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0, // pe_c2_r6::ConstVal
		1'bx, // pe_c2_r6::RegBConfig
		1'bx, // pe_c2_r6::RegAConfig
		1'bx, // pe_c2_r6::Reg7config
		1'bx, // pe_c2_r6::Reg6config
		1'bx, // pe_c2_r6::Reg5config
		1'bx, // pe_c2_r6::Reg4config
		1'bx, // pe_c2_r6::Reg3config
		1'bx, // pe_c2_r6::Reg2config
		1'bx, // pe_c2_r6::Reg1config
		1'bx, // pe_c2_r6::Reg0config
		1'bx, // pe_c2_r6::RESConfig
		1'b0, // pe_c2_r6::Mux7config
		1'bx, // pe_c2_r6::Mux6config
		1'bx, // pe_c2_r6::Mux5config
		1'bx, // pe_c2_r6::Mux4config
		1'bx, // pe_c2_r6::Mux3config
		1'bx, // pe_c2_r6::Mux2config
		1'bx, // pe_c2_r6::Mux1config
		1'bx, // pe_c2_r6::Mux0config
		1'bx,1'bx,1'bx,1'bx, // pe_c2_r6::ALUconfig
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux9config
		1'b1,1'b1,1'b0,1'b0, // crossbar::Mux8config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux7config
		1'b1,1'b0,1'b1,1'b0, // crossbar::Mux6config
		1'b0,1'b0,1'b0,1'b1, // crossbar::Mux5config
		1'b0,1'b1,1'b1,1'b0, // crossbar::Mux4config
		1'b1,1'b0,1'b0,1'b0, // crossbar::Mux3config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux2config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux1config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux0config
		1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0, // pe_c2_r5::ConstVal
		1'b1, // pe_c2_r5::RegBConfig
		1'bx, // pe_c2_r5::RegAConfig
		1'bx, // pe_c2_r5::Reg7config
		1'bx, // pe_c2_r5::Reg6config
		1'bx, // pe_c2_r5::Reg5config
		1'bx, // pe_c2_r5::Reg4config
		1'bx, // pe_c2_r5::Reg3config
		1'bx, // pe_c2_r5::Reg2config
		1'bx, // pe_c2_r5::Reg1config
		1'bx, // pe_c2_r5::Reg0config
		1'bx, // pe_c2_r5::RESConfig
		1'bx, // pe_c2_r5::Mux7config
		1'b0, // pe_c2_r5::Mux6config
		1'b0, // pe_c2_r5::Mux5config
		1'bx, // pe_c2_r5::Mux4config
		1'b0, // pe_c2_r5::Mux3config
		1'bx, // pe_c2_r5::Mux2config
		1'b0, // pe_c2_r5::Mux1config
		1'bx, // pe_c2_r5::Mux0config
		1'b0,1'b0,1'b1,1'b1, // pe_c2_r5::ALUconfig
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux9config
		1'b0,1'b0,1'b1,1'b0, // crossbar::Mux8config
		1'b1,1'b0,1'b1,1'b0, // crossbar::Mux7config
		1'b0,1'b0,1'b0,1'b0, // crossbar::Mux6config
		1'b1,1'b0,1'b0,1'b1, // crossbar::Mux5config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux4config
		1'b1,1'b0,1'b0,1'b0, // crossbar::Mux3config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux2config
		1'b1,1'b0,1'b0,1'b1, // crossbar::Mux1config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux0config
		1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0, // pe_c2_r4::ConstVal
		1'b1, // pe_c2_r4::RegBConfig
		1'bx, // pe_c2_r4::RegAConfig
		1'bx, // pe_c2_r4::Reg7config
		1'bx, // pe_c2_r4::Reg6config
		1'bx, // pe_c2_r4::Reg5config
		1'bx, // pe_c2_r4::Reg4config
		1'bx, // pe_c2_r4::Reg3config
		1'bx, // pe_c2_r4::Reg2config
		1'b1, // pe_c2_r4::Reg1config
		1'b1, // pe_c2_r4::Reg0config
		1'b1, // pe_c2_r4::RESConfig
		1'bx, // pe_c2_r4::Mux7config
		1'bx, // pe_c2_r4::Mux6config
		1'b0, // pe_c2_r4::Mux5config
		1'b0, // pe_c2_r4::Mux4config
		1'bx, // pe_c2_r4::Mux3config
		1'bx, // pe_c2_r4::Mux2config
		1'b1, // pe_c2_r4::Mux1config
		1'b1, // pe_c2_r4::Mux0config
		1'b0,1'b0,1'b1,1'b1, // pe_c2_r4::ALUconfig
		1'b1,1'b0,1'b1,1'b0, // crossbar::Mux9config
		1'b0,1'b0,1'b0,1'b0, // crossbar::Mux8config
		1'b0,1'b0,1'b1,1'b0, // crossbar::Mux7config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux6config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux5config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux4config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux3config
		1'b1,1'b0,1'b0,1'b1, // crossbar::Mux2config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux1config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux0config
		1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0, // pe_c2_r3::ConstVal
		1'b1, // pe_c2_r3::RegBConfig
		1'b1, // pe_c2_r3::RegAConfig
		1'bx, // pe_c2_r3::Reg7config
		1'bx, // pe_c2_r3::Reg6config
		1'bx, // pe_c2_r3::Reg5config
		1'bx, // pe_c2_r3::Reg4config
		1'bx, // pe_c2_r3::Reg3config
		1'bx, // pe_c2_r3::Reg2config
		1'bx, // pe_c2_r3::Reg1config
		1'bx, // pe_c2_r3::Reg0config
		1'b1, // pe_c2_r3::RESConfig
		1'bx, // pe_c2_r3::Mux7config
		1'bx, // pe_c2_r3::Mux6config
		1'b0, // pe_c2_r3::Mux5config
		1'b0, // pe_c2_r3::Mux4config
		1'bx, // pe_c2_r3::Mux3config
		1'bx, // pe_c2_r3::Mux2config
		1'bx, // pe_c2_r3::Mux1config
		1'b0, // pe_c2_r3::Mux0config
		1'b0,1'b0,1'b0,1'b0, // pe_c2_r3::ALUconfig
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux9config
		1'b1,1'b1,1'b0,1'b0, // crossbar::Mux8config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux7config
		1'b1,1'b0,1'b0,1'b1, // crossbar::Mux6config
		1'b1,1'b0,1'b0,1'b1, // crossbar::Mux5config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux4config
		1'b1,1'b0,1'b1,1'b0, // crossbar::Mux3config
		1'b0,1'b0,1'b1,1'b0, // crossbar::Mux2config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux1config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux0config
		1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0, // pe_c2_r2::ConstVal
		1'b1, // pe_c2_r2::RegBConfig
		1'bx, // pe_c2_r2::RegAConfig
		1'bx, // pe_c2_r2::Reg7config
		1'bx, // pe_c2_r2::Reg6config
		1'bx, // pe_c2_r2::Reg5config
		1'b1, // pe_c2_r2::Reg4config
		1'bx, // pe_c2_r2::Reg3config
		1'bx, // pe_c2_r2::Reg2config
		1'bx, // pe_c2_r2::Reg1config
		1'bx, // pe_c2_r2::Reg0config
		1'b1, // pe_c2_r2::RESConfig
		1'bx, // pe_c2_r2::Mux7config
		1'bx, // pe_c2_r2::Mux6config
		1'b0, // pe_c2_r2::Mux5config
		1'b1, // pe_c2_r2::Mux4config
		1'b0, // pe_c2_r2::Mux3config
		1'bx, // pe_c2_r2::Mux2config
		1'bx, // pe_c2_r2::Mux1config
		1'bx, // pe_c2_r2::Mux0config
		1'b1,1'b1,1'b0,1'b1, // pe_c2_r2::ALUconfig
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux9config
		1'b1,1'b1,1'b0,1'b0, // crossbar::Mux8config
		1'b1,1'b0,1'b0,1'b0, // crossbar::Mux7config
		1'b0,1'b0,1'b0,1'b1, // crossbar::Mux6config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux5config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux4config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux3config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux2config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux1config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux0config
		1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0, // pe_c2_r1::ConstVal
		1'b1, // pe_c2_r1::RegBConfig
		1'bx, // pe_c2_r1::RegAConfig
		1'bx, // pe_c2_r1::Reg7config
		1'bx, // pe_c2_r1::Reg6config
		1'bx, // pe_c2_r1::Reg5config
		1'bx, // pe_c2_r1::Reg4config
		1'bx, // pe_c2_r1::Reg3config
		1'bx, // pe_c2_r1::Reg2config
		1'bx, // pe_c2_r1::Reg1config
		1'bx, // pe_c2_r1::Reg0config
		1'bx, // pe_c2_r1::RESConfig
		1'bx, // pe_c2_r1::Mux7config
		1'bx, // pe_c2_r1::Mux6config
		1'bx, // pe_c2_r1::Mux5config
		1'bx, // pe_c2_r1::Mux4config
		1'b0, // pe_c2_r1::Mux3config
		1'bx, // pe_c2_r1::Mux2config
		1'b0, // pe_c2_r1::Mux1config
		1'bx, // pe_c2_r1::Mux0config
		1'b1,1'b1,1'b0,1'b1, // pe_c2_r1::ALUconfig
		1'b0,1'b0,1'b1,1'b0, // crossbar::Mux7config
		1'b1,1'b1,1'b0,1'b0, // crossbar::Mux6config
		1'b1,1'b0,1'b0,1'b0, // crossbar::Mux5config
		1'b1,1'b0,1'b1,1'b0, // crossbar::Mux4config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux3config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux2config
		1'b0,1'b1,1'b1,1'b0, // crossbar::Mux1config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux0config
		1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0, // pe_c2_r0::ConstVal
		1'b1, // pe_c2_r0::RegBConfig
		1'b1, // pe_c2_r0::RegAConfig
		1'b1, // pe_c2_r0::Reg7config
		1'bx, // pe_c2_r0::Reg6config
		1'b1, // pe_c2_r0::Reg3config
		1'bx, // pe_c2_r0::Reg2config
		1'bx, // pe_c2_r0::Reg1config
		1'bx, // pe_c2_r0::Reg0config
		1'bx, // pe_c2_r0::RESConfig
		1'b1, // pe_c2_r0::Mux7config
		1'b0, // pe_c2_r0::Mux6config
		1'b1, // pe_c2_r0::Mux3config
		1'bx, // pe_c2_r0::Mux2config
		1'b0, // pe_c2_r0::Mux1config
		1'bx, // pe_c2_r0::Mux0config
		1'b1,1'b0,1'b0,1'b0, // pe_c2_r0::ALUconfig
		1'b0,1'b0,1'b0,1'b0, // crossbar::Mux7config
		1'b1,1'b0,1'b0,1'b0, // crossbar::Mux6config
		1'b1,1'b1,1'b0,1'b0, // crossbar::Mux5config
		1'b1,1'b1,1'b1,1'b0, // crossbar::Mux4config
		1'b0,1'b1,1'b0,1'b0, // crossbar::Mux3config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux2config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux1config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux0config
		1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0, // pe_c1_r7::ConstVal
		1'b1, // pe_c1_r7::RegBConfig
		1'b1, // pe_c1_r7::RegAConfig
		1'bx, // pe_c1_r7::Reg5config
		1'bx, // pe_c1_r7::Reg4config
		1'bx, // pe_c1_r7::Reg3config
		1'b1, // pe_c1_r7::Reg2config
		1'bx, // pe_c1_r7::Reg1config
		1'bx, // pe_c1_r7::Reg0config
		1'b1, // pe_c1_r7::RESConfig
		1'bx, // pe_c1_r7::Mux5config
		1'bx, // pe_c1_r7::Mux4config
		1'b0, // pe_c1_r7::Mux3config
		1'b1, // pe_c1_r7::Mux2config
		1'b0, // pe_c1_r7::Mux1config
		1'b0, // pe_c1_r7::Mux0config
		1'b0,1'b1,1'b0,1'b1, // pe_c1_r7::ALUconfig
		1'b0,1'b1,1'b1,1'b0, // crossbar::Mux9config
		1'b0,1'b0,1'b0,1'b1, // crossbar::Mux8config
		1'b1,1'b0,1'b0,1'b1, // crossbar::Mux7config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux6config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux5config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux4config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux3config
		1'b1,1'b0,1'b0,1'b1, // crossbar::Mux2config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux1config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux0config
		1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0, // pe_c1_r6::ConstVal
		1'b1, // pe_c1_r6::RegBConfig
		1'b1, // pe_c1_r6::RegAConfig
		1'bx, // pe_c1_r6::Reg7config
		1'bx, // pe_c1_r6::Reg6config
		1'bx, // pe_c1_r6::Reg5config
		1'bx, // pe_c1_r6::Reg4config
		1'bx, // pe_c1_r6::Reg3config
		1'bx, // pe_c1_r6::Reg2config
		1'bx, // pe_c1_r6::Reg1config
		1'bx, // pe_c1_r6::Reg0config
		1'b1, // pe_c1_r6::RESConfig
		1'bx, // pe_c1_r6::Mux7config
		1'b0, // pe_c1_r6::Mux6config
		1'bx, // pe_c1_r6::Mux5config
		1'bx, // pe_c1_r6::Mux4config
		1'bx, // pe_c1_r6::Mux3config
		1'bx, // pe_c1_r6::Mux2config
		1'bx, // pe_c1_r6::Mux1config
		1'bx, // pe_c1_r6::Mux0config
		1'b0,1'b0,1'b0,1'b0, // pe_c1_r6::ALUconfig
		1'b1,1'b0,1'b0,1'b0, // crossbar::Mux9config
		1'b0,1'b0,1'b0,1'b0, // crossbar::Mux8config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux7config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux6config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux5config
		1'b0,1'b0,1'b0,1'b1, // crossbar::Mux4config
		1'b1,1'b0,1'b1,1'b0, // crossbar::Mux3config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux2config
		1'b0,1'b0,1'b1,1'b0, // crossbar::Mux1config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux0config
		1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0, // pe_c1_r5::ConstVal
		1'b1, // pe_c1_r5::RegBConfig
		1'b1, // pe_c1_r5::RegAConfig
		1'bx, // pe_c1_r5::Reg7config
		1'bx, // pe_c1_r5::Reg6config
		1'bx, // pe_c1_r5::Reg5config
		1'bx, // pe_c1_r5::Reg4config
		1'bx, // pe_c1_r5::Reg3config
		1'bx, // pe_c1_r5::Reg2config
		1'bx, // pe_c1_r5::Reg1config
		1'b1, // pe_c1_r5::Reg0config
		1'bx, // pe_c1_r5::RESConfig
		1'bx, // pe_c1_r5::Mux7config
		1'bx, // pe_c1_r5::Mux6config
		1'b0, // pe_c1_r5::Mux5config
		1'b0, // pe_c1_r5::Mux4config
		1'bx, // pe_c1_r5::Mux3config
		1'bx, // pe_c1_r5::Mux2config
		1'b0, // pe_c1_r5::Mux1config
		1'b1, // pe_c1_r5::Mux0config
		1'b1,1'b0,1'b1,1'b1, // pe_c1_r5::ALUconfig
		1'b0,1'b1,1'b1,1'b0, // crossbar::Mux9config
		1'b0,1'b0,1'b0,1'b0, // crossbar::Mux8config
		1'b1,1'b0,1'b1,1'b0, // crossbar::Mux7config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux6config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux5config
		1'b1,1'b0,1'b0,1'b0, // crossbar::Mux4config
		1'b0,1'b1,1'b1,1'b0, // crossbar::Mux3config
		1'b0,1'b0,1'b1,1'b0, // crossbar::Mux2config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux1config
		1'b1,1'b0,1'b0,1'b1, // crossbar::Mux0config
		1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0, // pe_c1_r4::ConstVal
		1'b1, // pe_c1_r4::RegBConfig
		1'b1, // pe_c1_r4::RegAConfig
		1'bx, // pe_c1_r4::Reg7config
		1'bx, // pe_c1_r4::Reg6config
		1'bx, // pe_c1_r4::Reg5config
		1'bx, // pe_c1_r4::Reg4config
		1'bx, // pe_c1_r4::Reg3config
		1'bx, // pe_c1_r4::Reg2config
		1'bx, // pe_c1_r4::Reg1config
		1'b1, // pe_c1_r4::Reg0config
		1'b1, // pe_c1_r4::RESConfig
		1'bx, // pe_c1_r4::Mux7config
		1'b0, // pe_c1_r4::Mux6config
		1'b0, // pe_c1_r4::Mux5config
		1'b0, // pe_c1_r4::Mux4config
		1'bx, // pe_c1_r4::Mux3config
		1'bx, // pe_c1_r4::Mux2config
		1'b0, // pe_c1_r4::Mux1config
		1'b1, // pe_c1_r4::Mux0config
		1'b0,1'b0,1'b0,1'b0, // pe_c1_r4::ALUconfig
		1'b0,1'b0,1'b0,1'b0, // crossbar::Mux9config
		1'b1,1'b1,1'b1,1'b0, // crossbar::Mux8config
		1'b0,1'b0,1'b1,1'b0, // crossbar::Mux7config
		1'b1,1'b1,1'b0,1'b0, // crossbar::Mux6config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux5config
		1'b0,1'b0,1'b0,1'b1, // crossbar::Mux4config
		1'b0,1'b1,1'b0,1'b0, // crossbar::Mux3config
		1'b0,1'b0,1'b1,1'b0, // crossbar::Mux2config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux1config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux0config
		1'b1,1'b1,1'b1,1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0, // pe_c1_r3::ConstVal
		1'b1, // pe_c1_r3::RegBConfig
		1'b1, // pe_c1_r3::RegAConfig
		1'bx, // pe_c1_r3::Reg7config
		1'bx, // pe_c1_r3::Reg6config
		1'bx, // pe_c1_r3::Reg5config
		1'bx, // pe_c1_r3::Reg4config
		1'bx, // pe_c1_r3::Reg3config
		1'bx, // pe_c1_r3::Reg2config
		1'bx, // pe_c1_r3::Reg1config
		1'bx, // pe_c1_r3::Reg0config
		1'bx, // pe_c1_r3::RESConfig
		1'b0, // pe_c1_r3::Mux7config
		1'bx, // pe_c1_r3::Mux6config
		1'bx, // pe_c1_r3::Mux5config
		1'b0, // pe_c1_r3::Mux4config
		1'b0, // pe_c1_r3::Mux3config
		1'b0, // pe_c1_r3::Mux2config
		1'bx, // pe_c1_r3::Mux1config
		1'b0, // pe_c1_r3::Mux0config
		1'b1,1'b0,1'b1,1'b1, // pe_c1_r3::ALUconfig
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux9config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux8config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux7config
		1'b0,1'b0,1'b1,1'b0, // crossbar::Mux6config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux5config
		1'b1,1'b0,1'b0,1'b0, // crossbar::Mux4config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux3config
		1'b1,1'b0,1'b1,1'b0, // crossbar::Mux2config
		1'b1,1'b1,1'b0,1'b0, // crossbar::Mux1config
		1'b0,1'b0,1'b1,1'b0, // crossbar::Mux0config
		1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0, // pe_c1_r2::ConstVal
		1'bx, // pe_c1_r2::RegBConfig
		1'bx, // pe_c1_r2::RegAConfig
		1'bx, // pe_c1_r2::Reg7config
		1'bx, // pe_c1_r2::Reg6config
		1'bx, // pe_c1_r2::Reg5config
		1'bx, // pe_c1_r2::Reg4config
		1'bx, // pe_c1_r2::Reg3config
		1'bx, // pe_c1_r2::Reg2config
		1'bx, // pe_c1_r2::Reg1config
		1'bx, // pe_c1_r2::Reg0config
		1'bx, // pe_c1_r2::RESConfig
		1'bx, // pe_c1_r2::Mux7config
		1'bx, // pe_c1_r2::Mux6config
		1'b0, // pe_c1_r2::Mux5config
		1'b0, // pe_c1_r2::Mux4config
		1'b0, // pe_c1_r2::Mux3config
		1'bx, // pe_c1_r2::Mux2config
		1'b0, // pe_c1_r2::Mux1config
		1'bx, // pe_c1_r2::Mux0config
		1'bx,1'bx,1'bx,1'bx, // pe_c1_r2::ALUconfig
		1'b0,1'b1,1'b0,1'b0, // crossbar::Mux9config
		1'b1,1'b0,1'b1,1'b0, // crossbar::Mux8config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux7config
		1'b0,1'b0,1'b1,1'b0, // crossbar::Mux6config
		1'b0,1'b1,1'b0,1'b1, // crossbar::Mux5config
		1'b0,1'b0,1'b0,1'b1, // crossbar::Mux4config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux3config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux2config
		1'b1,1'b1,1'b1,1'b0, // crossbar::Mux1config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux0config
		1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0, // pe_c1_r1::ConstVal
		1'b1, // pe_c1_r1::RegBConfig
		1'b1, // pe_c1_r1::RegAConfig
		1'bx, // pe_c1_r1::Reg7config
		1'bx, // pe_c1_r1::Reg6config
		1'bx, // pe_c1_r1::Reg5config
		1'bx, // pe_c1_r1::Reg4config
		1'bx, // pe_c1_r1::Reg3config
		1'b1, // pe_c1_r1::Reg2config
		1'bx, // pe_c1_r1::Reg1config
		1'bx, // pe_c1_r1::Reg0config
		1'bx, // pe_c1_r1::RESConfig
		1'b0, // pe_c1_r1::Mux7config
		1'bx, // pe_c1_r1::Mux6config
		1'b0, // pe_c1_r1::Mux5config
		1'b0, // pe_c1_r1::Mux4config
		1'bx, // pe_c1_r1::Mux3config
		1'b1, // pe_c1_r1::Mux2config
		1'bx, // pe_c1_r1::Mux1config
		1'bx, // pe_c1_r1::Mux0config
		1'b0,1'b1,1'b0,1'b1, // pe_c1_r1::ALUconfig
		1'b1,1'b0,1'b1,1'b0, // crossbar::Mux7config
		1'b0,1'b0,1'b0,1'b0, // crossbar::Mux6config
		1'b1,1'b1,1'b1,1'b0, // crossbar::Mux5config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux4config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux3config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux2config
		1'b1,1'b1,1'b0,1'b0, // crossbar::Mux1config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux0config
		1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0, // pe_c1_r0::ConstVal
		1'b1, // pe_c1_r0::RegBConfig
		1'b1, // pe_c1_r0::RegAConfig
		1'b1, // pe_c1_r0::Reg7config
		1'bx, // pe_c1_r0::Reg6config
		1'bx, // pe_c1_r0::Reg3config
		1'bx, // pe_c1_r0::Reg2config
		1'bx, // pe_c1_r0::Reg1config
		1'bx, // pe_c1_r0::Reg0config
		1'b1, // pe_c1_r0::RESConfig
		1'b1, // pe_c1_r0::Mux7config
		1'bx, // pe_c1_r0::Mux6config
		1'b0, // pe_c1_r0::Mux3config
		1'bx, // pe_c1_r0::Mux2config
		1'bx, // pe_c1_r0::Mux1config
		1'b0, // pe_c1_r0::Mux0config
		1'b0,1'b1,1'b0,1'b1, // pe_c1_r0::ALUconfig
		1'b0,1'b0,1'b1, // crossbar::Mux6config
		1'b1,1'b0,1'b0, // crossbar::Mux5config
		1'bx,1'bx,1'bx, // crossbar::Mux4config
		1'b0,1'b1,1'b1, // crossbar::Mux3config
		1'bx,1'bx,1'bx, // crossbar::Mux2config
		1'b1,1'b1,1'b1, // crossbar::Mux1config
		1'b0,1'b1,1'b0, // crossbar::Mux0config
		1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0, // pe_c0_r7::ConstVal
		1'b1, // pe_c0_r7::RegBConfig
		1'b1, // pe_c0_r7::RegAConfig
		1'bx, // pe_c0_r7::Reg5config
		1'bx, // pe_c0_r7::Reg3config
		1'bx, // pe_c0_r7::Reg2config
		1'b1, // pe_c0_r7::Reg1config
		1'bx, // pe_c0_r7::Reg0config
		1'b1, // pe_c0_r7::RESConfig
		1'b0, // pe_c0_r7::Mux5config
		1'bx, // pe_c0_r7::Mux3config
		1'b0, // pe_c0_r7::Mux2config
		1'b1, // pe_c0_r7::Mux1config
		1'bx, // pe_c0_r7::Mux0config
		1'b0,1'b1,1'b0,1'b1, // pe_c0_r7::ALUconfig
		1'b0,1'b0,1'b0,1'b0, // crossbar::Mux7config
		1'b0,1'b1,1'b0,1'b0, // crossbar::Mux6config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux5config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux4config
		1'b1,1'b0,1'b1,1'b0, // crossbar::Mux3config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux2config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux1config
		1'b0,1'b1,1'b1,1'b0, // crossbar::Mux0config
		1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0, // pe_c0_r6::ConstVal
		1'b1, // pe_c0_r6::RegBConfig
		1'b1, // pe_c0_r6::RegAConfig
		1'b1, // pe_c0_r6::Reg6config
		1'bx, // pe_c0_r6::Reg5config
		1'bx, // pe_c0_r6::Reg3config
		1'b1, // pe_c0_r6::Reg2config
		1'bx, // pe_c0_r6::Reg1config
		1'bx, // pe_c0_r6::Reg0config
		1'bx, // pe_c0_r6::RESConfig
		1'b1, // pe_c0_r6::Mux6config
		1'bx, // pe_c0_r6::Mux5config
		1'bx, // pe_c0_r6::Mux3config
		1'b1, // pe_c0_r6::Mux2config
		1'bx, // pe_c0_r6::Mux1config
		1'b0, // pe_c0_r6::Mux0config
		1'b0,1'b1,1'b0,1'b1, // pe_c0_r6::ALUconfig
		1'b1,1'b0,1'b0,1'b0, // crossbar::Mux7config
		1'b0,1'b0,1'b0,1'b0, // crossbar::Mux6config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux5config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux4config
		1'b0,1'b1,1'b0,1'b0, // crossbar::Mux3config
		1'b0,1'b0,1'b1,1'b0, // crossbar::Mux2config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux1config
		1'b0,1'b1,1'b1,1'b0, // crossbar::Mux0config
		1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0, // pe_c0_r5::ConstVal
		1'b1, // pe_c0_r5::RegBConfig
		1'b1, // pe_c0_r5::RegAConfig
		1'bx, // pe_c0_r5::Reg6config
		1'bx, // pe_c0_r5::Reg5config
		1'bx, // pe_c0_r5::Reg3config
		1'bx, // pe_c0_r5::Reg2config
		1'bx, // pe_c0_r5::Reg1config
		1'b1, // pe_c0_r5::Reg0config
		1'bx, // pe_c0_r5::RESConfig
		1'bx, // pe_c0_r5::Mux6config
		1'b0, // pe_c0_r5::Mux5config
		1'bx, // pe_c0_r5::Mux3config
		1'b0, // pe_c0_r5::Mux2config
		1'b0, // pe_c0_r5::Mux1config
		1'b1, // pe_c0_r5::Mux0config
		1'b0,1'b0,1'b0,1'b1, // pe_c0_r5::ALUconfig
		1'b1,1'b0,1'b0,1'b0, // crossbar::Mux7config
		1'b0,1'b0,1'b1,1'b0, // crossbar::Mux6config
		1'b0,1'b0,1'b0,1'b0, // crossbar::Mux5config
		1'b0,1'b1,1'b0,1'b0, // crossbar::Mux4config
		1'b1,1'b0,1'b1,1'b0, // crossbar::Mux3config
		1'b1,1'b1,1'b1,1'b0, // crossbar::Mux2config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux1config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux0config
		1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0, // pe_c0_r4::ConstVal
		1'b1, // pe_c0_r4::RegBConfig
		1'b1, // pe_c0_r4::RegAConfig
		1'bx, // pe_c0_r4::Reg6config
		1'b1, // pe_c0_r4::Reg5config
		1'bx, // pe_c0_r4::Reg3config
		1'bx, // pe_c0_r4::Reg2config
		1'bx, // pe_c0_r4::Reg1config
		1'bx, // pe_c0_r4::Reg0config
		1'b1, // pe_c0_r4::RESConfig
		1'b0, // pe_c0_r4::Mux6config
		1'b1, // pe_c0_r4::Mux5config
		1'bx, // pe_c0_r4::Mux3config
		1'b0, // pe_c0_r4::Mux2config
		1'b0, // pe_c0_r4::Mux1config
		1'b0, // pe_c0_r4::Mux0config
		1'b1,1'b0,1'b0,1'b0, // pe_c0_r4::ALUconfig
		1'b1,1'b0,1'b1,1'b0, // crossbar::Mux7config
		1'b1,1'b0,1'b0,1'b0, // crossbar::Mux6config
		1'b1,1'b1,1'b1,1'b0, // crossbar::Mux5config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux4config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux3config
		1'b1,1'b1,1'b0,1'b0, // crossbar::Mux2config
		1'b0,1'b0,1'b0,1'b0, // crossbar::Mux1config
		1'b1,1'b1,1'b0,1'b0, // crossbar::Mux0config
		1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0, // pe_c0_r3::ConstVal
		1'b1, // pe_c0_r3::RegBConfig
		1'b1, // pe_c0_r3::RegAConfig
		1'bx, // pe_c0_r3::Reg6config
		1'bx, // pe_c0_r3::Reg5config
		1'bx, // pe_c0_r3::Reg3config
		1'bx, // pe_c0_r3::Reg2config
		1'bx, // pe_c0_r3::Reg1config
		1'bx, // pe_c0_r3::Reg0config
		1'b1, // pe_c0_r3::RESConfig
		1'b0, // pe_c0_r3::Mux6config
		1'bx, // pe_c0_r3::Mux5config
		1'b0, // pe_c0_r3::Mux3config
		1'bx, // pe_c0_r3::Mux2config
		1'b0, // pe_c0_r3::Mux1config
		1'b0, // pe_c0_r3::Mux0config
		1'b0,1'b0,1'b0,1'b1, // pe_c0_r3::ALUconfig
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux7config
		1'b0,1'b0,1'b0,1'b0, // crossbar::Mux6config
		1'b0,1'b1,1'b1,1'b0, // crossbar::Mux5config
		1'b0,1'b1,1'b0,1'b0, // crossbar::Mux4config
		1'b1,1'b0,1'b1,1'b0, // crossbar::Mux3config
		1'b1,1'b1,1'b0,1'b0, // crossbar::Mux2config
		1'b1,1'b1,1'b0,1'b0, // crossbar::Mux1config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux0config
		1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0, // pe_c0_r2::ConstVal
		1'b1, // pe_c0_r2::RegBConfig
		1'bx, // pe_c0_r2::RegAConfig
		1'bx, // pe_c0_r2::Reg6config
		1'bx, // pe_c0_r2::Reg5config
		1'bx, // pe_c0_r2::Reg3config
		1'bx, // pe_c0_r2::Reg2config
		1'bx, // pe_c0_r2::Reg1config
		1'b1, // pe_c0_r2::Reg0config
		1'bx, // pe_c0_r2::RESConfig
		1'b0, // pe_c0_r2::Mux6config
		1'bx, // pe_c0_r2::Mux5config
		1'b0, // pe_c0_r2::Mux3config
		1'b0, // pe_c0_r2::Mux2config
		1'bx, // pe_c0_r2::Mux1config
		1'b1, // pe_c0_r2::Mux0config
		1'b1,1'b1,1'b0,1'b1, // pe_c0_r2::ALUconfig
		1'b1,1'b0,1'b1,1'b0, // crossbar::Mux7config
		1'b0,1'b1,1'b1,1'b0, // crossbar::Mux6config
		1'b0,1'b1,1'b1,1'b0, // crossbar::Mux5config
		1'b1,1'b1,1'b1,1'b0, // crossbar::Mux4config
		1'b0,1'b0,1'b1,1'b0, // crossbar::Mux3config
		1'b1,1'b1,1'b0,1'b0, // crossbar::Mux2config
		1'bx,1'bx,1'bx,1'bx, // crossbar::Mux1config
		1'b1,1'b1,1'b0,1'b0, // crossbar::Mux0config
		1'b1,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0, // pe_c0_r1::ConstVal
		1'b1, // pe_c0_r1::RegBConfig
		1'b1, // pe_c0_r1::RegAConfig
		1'bx, // pe_c0_r1::Reg6config
		1'bx, // pe_c0_r1::Reg5config
		1'b1, // pe_c0_r1::Reg3config
		1'bx, // pe_c0_r1::Reg2config
		1'bx, // pe_c0_r1::Reg1config
		1'bx, // pe_c0_r1::Reg0config
		1'b1, // pe_c0_r1::RESConfig
		1'b0, // pe_c0_r1::Mux6config
		1'b0, // pe_c0_r1::Mux5config
		1'b1, // pe_c0_r1::Mux3config
		1'bx, // pe_c0_r1::Mux2config
		1'bx, // pe_c0_r1::Mux1config
		1'bx, // pe_c0_r1::Mux0config
		1'b0,1'b0,1'b0,1'b0, // pe_c0_r1::ALUconfig
		1'bx,1'bx,1'bx, // crossbar::Mux6config
		1'b0,1'b1,1'b0, // crossbar::Mux5config
		1'b1,1'b0,1'b1, // crossbar::Mux4config
		1'b0,1'b0,1'b1, // crossbar::Mux3config
		1'bx,1'bx,1'bx, // crossbar::Mux2config
		1'b0,1'b1,1'b1, // crossbar::Mux1config
		1'bx,1'bx,1'bx, // crossbar::Mux0config
		1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0, // pe_c0_r0::ConstVal
		1'b1, // pe_c0_r0::RegBConfig
		1'bx, // pe_c0_r0::RegAConfig
		1'bx, // pe_c0_r0::Reg6config
		1'bx, // pe_c0_r0::Reg3config
		1'b1, // pe_c0_r0::Reg2config
		1'bx, // pe_c0_r0::Reg1config
		1'bx, // pe_c0_r0::Reg0config
		1'b1, // pe_c0_r0::RESConfig
		1'b0, // pe_c0_r0::Mux6config
		1'bx, // pe_c0_r0::Mux3config
		1'b1, // pe_c0_r0::Mux2config
		1'bx, // pe_c0_r0::Mux1config
		1'bx, // pe_c0_r0::Mux0config
		1'b0,1'b0,1'b1,1'b1, // pe_c0_r0::ALUconfig
		1'b0, // mem_7::WriteRq
		1'bx,1'bx,1'bx, // mem_7::MuxData
		1'bx,1'bx,1'bx, // mem_7::MuxAddr
		1'b0, // mem_6::WriteRq
		1'bx,1'bx,1'bx, // mem_6::MuxData
		1'bx,1'bx,1'bx, // mem_6::MuxAddr
		1'b1, // mem_5::WriteRq
		1'b0,1'b1,1'b0, // mem_5::MuxData
		1'b1,1'b1,1'b1, // mem_5::MuxAddr
		1'b1, // mem_4::WriteRq
		1'b0,1'b0,1'b1, // mem_4::MuxData
		1'b0,1'b1,1'b1, // mem_4::MuxAddr
		1'b0, // mem_3::WriteRq
		1'bx,1'bx,1'bx, // mem_3::MuxData
		1'b0,1'b0,1'b0, // mem_3::MuxAddr
		1'b0, // mem_2::WriteRq
		1'bx,1'bx,1'bx, // mem_2::MuxData
		1'b1,1'b0,1'b1, // mem_2::MuxAddr
		1'b0, // mem_1::WriteRq
		1'bx,1'bx,1'bx, // mem_1::MuxData
		1'b1,1'b0,1'b0, // mem_1::MuxAddr
		1'b0, // mem_0::WriteRq
		1'bx,1'bx,1'bx, // mem_0::MuxData
		1'bx,1'bx,1'bx, // mem_0::MuxAddr
		1'bx, // io_top_7::RegOutConfig
		1'bx, // io_top_7::RegInConfig
		1'b0, // io_top_7::IOPinConfig
		1'bx, // io_top_6::RegOutConfig
		1'bx, // io_top_6::RegInConfig
		1'b0, // io_top_6::IOPinConfig
		1'bx, // io_top_5::RegOutConfig
		1'bx, // io_top_5::RegInConfig
		1'b0, // io_top_5::IOPinConfig
		1'bx, // io_top_4::RegOutConfig
		1'bx, // io_top_4::RegInConfig
		1'b0, // io_top_4::IOPinConfig
		1'b1, // io_top_3::RegOutConfig
		1'bx, // io_top_3::RegInConfig
		1'b0, // io_top_3::IOPinConfig
		1'bx, // io_top_2::RegOutConfig
		1'bx, // io_top_2::RegInConfig
		1'b0, // io_top_2::IOPinConfig
		1'b1, // io_top_1::RegOutConfig
		1'bx, // io_top_1::RegInConfig
		1'b0, // io_top_1::IOPinConfig
		1'bx, // io_top_0::RegOutConfig
		1'bx, // io_top_0::RegInConfig
		1'b0, // io_top_0::IOPinConfig
		1'bx, // io_right_7::RegOutConfig
		1'bx, // io_right_7::RegInConfig
		1'b0, // io_right_7::IOPinConfig
		1'bx, // io_right_6::RegOutConfig
		1'bx, // io_right_6::RegInConfig
		1'b0, // io_right_6::IOPinConfig
		1'bx, // io_right_5::RegOutConfig
		1'bx, // io_right_5::RegInConfig
		1'b0, // io_right_5::IOPinConfig
		1'bx, // io_right_4::RegOutConfig
		1'bx, // io_right_4::RegInConfig
		1'b0, // io_right_4::IOPinConfig
		1'bx, // io_right_3::RegOutConfig
		1'bx, // io_right_3::RegInConfig
		1'b0, // io_right_3::IOPinConfig
		1'bx, // io_right_2::RegOutConfig
		1'bx, // io_right_2::RegInConfig
		1'b0, // io_right_2::IOPinConfig
		1'bx, // io_right_1::RegOutConfig
		1'bx, // io_right_1::RegInConfig
		1'b0, // io_right_1::IOPinConfig
		1'bx, // io_right_0::RegOutConfig
		1'bx, // io_right_0::RegInConfig
		1'b0, // io_right_0::IOPinConfig
		1'bx, // io_bottom_7::RegOutConfig
		1'bx, // io_bottom_7::RegInConfig
		1'b0, // io_bottom_7::IOPinConfig
		1'bx, // io_bottom_6::RegOutConfig
		1'bx, // io_bottom_6::RegInConfig
		1'b0, // io_bottom_6::IOPinConfig
		1'bx, // io_bottom_5::RegOutConfig
		1'bx, // io_bottom_5::RegInConfig
		1'b0, // io_bottom_5::IOPinConfig
		1'bx, // io_bottom_4::RegOutConfig
		1'bx, // io_bottom_4::RegInConfig
		1'b0, // io_bottom_4::IOPinConfig
		1'b1, // io_bottom_3::RegOutConfig
		1'bx, // io_bottom_3::RegInConfig
		1'b0, // io_bottom_3::IOPinConfig
		1'bx, // io_bottom_2::RegOutConfig
		1'bx, // io_bottom_2::RegInConfig
		1'b0, // io_bottom_2::IOPinConfig
		1'b1, // io_bottom_1::RegOutConfig
		1'bx, // io_bottom_1::RegInConfig
		1'b0, // io_bottom_1::IOPinConfig
		1'b1, // io_bottom_0::RegOutConfig
		1'bx, // io_bottom_0::RegInConfig
		1'b0 // io_bottom_0::IOPinConfig
	};

	reg [31:0] next_pos;
	always @(posedge clock) begin
		if (sync_reset) begin
			next_pos <= 0;
			bitstream <= 1'b0;
			done <= 0;
		end else if (next_pos >= TOTAL_NUM_BITS) begin
			done <= 1;
			bitstream <= 1'b0;
		end else if (enable) begin
			bitstream <= storage[next_pos];
			next_pos <= next_pos + 1;
		end
	end
endmodule
